`timescale 1ns / 1ps

module tb_SpMV_ops();

	reg			i_clk;
	reg			i_rstn;
	reg         i_start;

	reg	[255:0]	i_read_data_A;
	reg [255:0]	i_read_data_B;

	wire [255:0] o_result;

	SpMV_ops uut(
		.i_clk(i_clk),
		.i_rstn(i_rstn),
		.i_start(i_start),
		
		.i_read_data_A(i_read_data_A),
		.i_read_data_B(i_read_data_B),

		.o_result(o_result)
	);

	initial begin
		i_clk = 1'b0; i_rstn = 1'b0; i_start = 1'b0;
		#30 i_rstn = 1'b1;
		#44 i_start = 1'b1;
	end

	always begin
		#5 i_clk = ~i_clk;
	end

	initial begin
		i_read_data_A = 0;
		i_read_data_B = 0;
		// A = Input Vector, B = Row Pointer
		#74   // A = [1, 3.1, 31, 0.41, 0.18, 6.31, 3, 8, 0, 1.2, 57.1, 31.3, 4.1, 1.2, 75, 31], B = [0, 0, 1, 2, 2, 2, 2, 3, 3, 3, 3, 4, 5, 5, 5, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
		i_read_data_A = 256'b0_10011_1111000000_0_10101_0010110000_0_01111_0011001101_0_10001_0000011010_0_10011_1111010011_0_10100_1100100011_0_01111_0011001101_0_00000_0000000000_0_10010_0000000000_0_10000_1000000000_0_10001_1001001111_0_01100_0111000011_0_01101_1010001111_0_10011_1111000000_0_10000_1000110011_0_01111_0000000000;
		i_read_data_B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000110_00000101_00000101_00000101_00000100_00000011_00000011_00000011_00000011_00000010_00000010_00000010_00000010_00000001_00000000_00000000;
		// A = Value, B = Column Index
		#15   // A = [1.03, 5.2, 7, 3.1, 10, 2], B = [ 0, 3, 7, 11, 14, 15]
		i_read_data_A = 256'b0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0_10000_0000000000_0_10010_0100000000_0_10000_1000110011_0_10001_1100000000_0_10001_0100110011_0_01111_0000011111;
		i_read_data_B = 256'b0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_1110_1101_1011_0111_0011_0000;
	end


//	initial begin
//		$dumpfile("tb_SpMV_ops.vcd");
//		$dumpvars(0,tb_SpMV_ops);
//	end


endmodule
