`timescale 1ns / 1ps

module tb_SpMV_ops_controller();

    reg i_clk;
    reg i_rstn;
    
    reg [255:0]             i_read_data_A;
    reg [255:0]             i_read_data_B;
    
    wire [4:0]              o_address_A;
    wire [4:0]              o_address_B;
    
    wire                    o_wr_en_A;
    wire                    o_wr_en_B;
    
    wire [2:0]              o_state;
    wire [3:0]              o_SRAM0_state;
    wire [3:0]              o_SRAM1_state;
    wire [3:0]              o_core_state;
    wire                    o_write_state;
    wire                    o_done;
   
   wire [255:0]             o_write_data_A;
   wire [255:0]             o_write_data_B;
   
   
   SpMV_ops_controller u0(
        .i_clk(i_clk),
        .i_rstn(i_rstn),
        .i_read_data_A(i_read_data_A),
        .i_read_data_B(i_read_data_B),
        .o_address_A(o_address_A),
        .o_address_B(o_address_B),
        .o_wr_en_A(o_wr_en_A),
        .o_wr_en_B(o_wr_en_B),
        .o_state(o_state),
        .o_SRAM0_state(o_SRAM0_state),
        .o_SRAM1_state(o_SRAM1_state),
        .o_core_state(o_core_state),
        .o_write_state(o_write_state),
        .o_done(o_done),
        .o_write_data_A(o_write_data_A),
        .o_write_data_B(o_write_data_B)
        );
 
     
     initial begin
        i_clk = 1'b0;
        i_rstn = 1'b0;
        #30
        i_rstn = 1'b1;
     end
 
     always begin
        #5 i_clk = ~i_clk;
     end

    initial begin
        i_read_data_A = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        i_read_data_B = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        
        // Polling DONE
        #103
        i_read_data_A = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001;
        
        #15
       i_read_data_A = 256'b0_10011_1111000000_0_10101_0010110000_0_01111_0011001101_0_10001_0000011010_0_10011_1111010011_0_10100_1100100011_0_01111_0011001101_0_00000_0000000000_0_10010_0000000000_0_10000_1000000000_0_10001_1001001111_0_01100_0111000011_0_01101_1010001111_0_10011_1111000000_0_10000_1000110011_0_01111_0000000000;
       i_read_data_B = 256'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000110_00000101_00000101_00000101_00000100_00000011_00000011_00000011_00000011_00000010_00000010_00000010_00000010_00000001_00000000_00000000;
        // A = Value, B = Column Index
        #10   // A = [1.03, 5.2, 7, 3.1, 10, 2], B = [ 0, 3, 7, 11, 14, 15]
        i_read_data_A = 256'b0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0_10000_0000000000_0_10010_0100000000_0_10000_1000110011_0_10001_1100000000_0_10001_0100110011_0_01111_0000011111;
        i_read_data_B = 256'b0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_1110_1101_1011_0111_0011_0000;
	end

  
endmodule
